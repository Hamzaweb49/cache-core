module tb_cache_controller;

    // TESTBENCH FOR CACHE CONTROLLER HERE

endmodule