module tb_ace_controller;

    // TESTBENCH FOR ACE CONTROLLER
endmodule