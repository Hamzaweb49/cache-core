module tb_cache_datapath;

    // TESTBENCH FOR DATAPATH HERE
endmodule