module tb_top_level;

    // TESTBENCH FOR TOP LEVEL HERE
endmodule